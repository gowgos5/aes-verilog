module AEScntx(
//from testbench
input  clk,
input  start,
input  rstn,
//to AEScore
output  accept,
output  [3:0] rndNo,
output  enbSB,
output  enbSR,
output  enbMC,
output  enbAR,
output  enbKS,
//to testbench
output  done,
output  [9:0] completed_round
);
////enter your code here
endmodule

module AddRndKey_top(
input  [127:0] ip,
input  [127:0] ip_key,
input  enable,
output  [127:0] op
);
////enter your code here
endmodule

module AESCore(
//from testbench
input  clk,
input  rstn,
input  [127:0] plain_text,
input  [127:0] cipher_key,
//from controller
input  accept,
input  [3:0] rndNo,
input  enbSB,
input  enbSR,
input  enbMC,
input  enbAR,
input  enbKS,
//to testbench
output [127:0] cipher_text
);
////enter your code here
endmodule

module AEScntx#(N=4)(
//from testbench
input bit clk,
input bit start,
input bit rstn,
//to AEScore
output bit accept,
output bit [3:0] rndNo,
output bit enbSB,
output bit enbSR,
output bit enbMC,
output bit enbAR,
output bit enbKS,
//to testbench
output bit done
);
////enter your code here
endmodule

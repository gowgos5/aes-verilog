module KeySchedule_top(
input  [127:0] ip_key,
input  enable,
input  [3:0] rndNo,
output  [127:0] op_key
);
////enter your code here
endmodule

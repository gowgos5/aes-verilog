module subBytes_top(
input [127:0] ip,
input enable,
output [127:0] op
);
////enter your code here
endmodule
